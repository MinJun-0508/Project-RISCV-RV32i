`timescale 1ns / 1ps

module instr_mem (
    input  logic [31:0] instr_rAddr,
    output logic [31:0] instr_code
);
    logic [31:0] rom[0:63];

    initial begin
        // 32'b imm(7bit) _ rs2(5bit) _ rs1(5bit) _ funct3(3bit) _ imm(5bit) _ opcode(7'b0100011)
        // R-type
        rom [0] = 32'b0000000_00010_00011_000_00001_0110011; //  add x1, x3, x2  | rd = 3 + 2  
        rom [1] = 32'b0100000_00010_00011_000_00001_0110011; //  sub x1, x3, x2  | rd = 3 - 2 
        rom [2] = 32'b0000000_00010_00011_001_00001_0110011; //  sll x1, x3, x2  | rd = 3 << 2  
        rom [3] = 32'b0000000_00010_00011_100_00001_0110011; //  xor x1, x3, x2  | rd = 3 ^ 2
        rom [4] = 32'b0000000_00010_00011_101_00001_0110011; //  srl x1, x3, x2  | rd = 3 >> 2
        rom [5] = 32'b0100000_00010_00011_101_00001_0110011; //  sra x1, x3, x2  | rd = 3 >> 2   
        rom [6] = 32'b0000000_00010_00011_110_00001_0110011; //  or  x1, x3, x2  | rd = 3 | 2   
        rom [7] = 32'b0000000_00010_00011_111_00001_0110011; //  and x1, x3, x2  | rd = 3 & 2  
        rom [8] = 32'b0000000_00010_00100_010_00001_0110011; //  slt x1, x4, x2  | rd = (-1 < 2) ? 1:0
        rom [9] = 32'b0000000_00010_00100_011_00001_0110011; // sltu x1, x4, x2  | rd = (2^32 - 1 < 2) ? 1:0


        // imm[7]_rs2[5]_rs1[5]_funct3[3]_imm[5]_opcode
        // S-type
        rom[0] = 32'b0000000_00010_00001_000_00001_0100011; // sb x8, 1(x1) | M[0+2][0:7]  = rs2[0:7]
        rom[1] = 32'b0000000_00010_00001_001_00001_0100011; // sh x8, 1(x1) | M[0+2][0:15] = rs2[0:15] 
        rom[2] = 32'b0000000_00010_00001_010_00001_0100011; // sw x8, 1(x1) | M[0+2][0:31] = rs2[0:31]

        //IL-type
        // rom [0] = 32'b000000000010_00000_000_00001_0000011; // lb  x1, 2(x0) | rd = M[0+2][0:7]
        // rom [1] = 32'b000000000010_00000_001_00001_0000011; // lh  x1, 2(x0) | rd = M[0+2][0:15]
        // rom [2] = 32'b000000000010_00000_010_00001_0000011; // lw  x1, 2(x0) | rd = M[0+2][0:31]
        // rom [3] = 32'b000000000010_00000_100_00001_0000011; // lbu x1, 2(x0) | rd = M[0+2][0:7]
        // rom [4] = 32'b000000000010_00000_101_00001_0000011; // lhu x1, 2(x0) | rd = M[0+2][0:15]

        // I-type, imm(12bit)_rs1(5bit)_funct3(3bit)_rd(5bit)_opcode(7bit)
        // I-type
        // rom[0] = 32'b000000001100_00110_000_00001_0010011; // addi  x1  x6  12 | rd = 6 + 12
        // rom[1] = 32'b111111111111_00110_010_00001_0010011; // slti  x1, x6, 12 | rd = (6 < -1)?1:0
        // rom[2] = 32'b111111111111_00110_011_00001_0010011; // sltiu x1, x6, 12 | rd = (6 < 2^32 - 1)?1:0
        // rom[3] = 32'b000000001100_00110_100_00001_0010011; // xori  x1, x6, 12 | rd = 6 ˆ 12
        // rom[4] = 32'b000000001100_00110_110_00001_0010011; // ori   x1, x6, 12 | rd = 6 | 12
        // rom[5] = 32'b000000001100_00110_111_00001_0010011; // andi  x1, x6, 12 | rd = 6 & 12
        // rom[6] = 32'b000000000001_00110_001_00001_0010011; // slli  x1, x6, 1  | rd = 6 << 1[0:4]
        // rom[7] = 32'b000000000010_00011_101_00010_0010011; // srli  x2, x3, 2  | rd = 3 >> 2[0:4]
        // rom[8] = 32'b010000000010_00011_101_00010_0010011; // srai  x2, x3, 2  | rd = 3 >> 2[0:4]

        // Branch
        // rom[0]  = 32'b0000000_00010_00010_000_10000_1100011;  //  beq x2, x2, 16 | if(2 == 2) PC += 16
        // rom[4]  = 32'b0000000_00010_00001_001_10000_1100011;  //  bne x1, x2, 16 | if(1 != 2) PC += 16
        // rom[8]  = 32'b0000000_00100_00010_100_10000_1100011;  //  blt x2, x4, 16 | if(2 <  4) PC += 16
        // rom[12] = 32'b0000000_00100_01000_101_10000_1100011;  //  bge x8, x4, 16 | if(8 >= 4) PC += 16
        // rom[16] = 32'b0000000_00100_00010_110_10000_1100011;  // bltu x2, x4, 16 | if(2 <  4) PC += 16
        // rom[20] = 32'b0000000_00010_00100_111_10000_1100011;  // bgeu x4, x2, 16 | if(4 >= 2) PC += 16


        // U-type
        // rom[0] = 32'b0000_0000_0000_0000_0001_00001_0110111; // lui   x1, 1 | rd = imm
        // rom[1] = 32'b0000_0000_0000_0000_0001_00001_0010111; // auipc x1, 1 | rd = PC + imm

        // jal, jarl
        rom[ 0] = 32'b0000_0010_0000_0000_0000_00001_1101111; // jal x1, 32      | rd = PC+4; PC += 32
        rom[ 8] = 32'b0000_0100_0000_00100_000_00001_1100111; // jalr x1, 64(x4) | rd = PC+4; PC = 4 + 64 
        rom[17] = 32'b0000000_00010_00011_000_00001_0110011;  // add x1, x3, x2  | rd = 3 + 2
    end

    assign instr_code = rom[instr_rAddr[31:2]];

endmodule
